module i2c_master (
	input CLOCK_50,
	inout SDA,
	output SCLs
);

endmodule